module A;
always @* begin
end
endmodule
