module A;
always_comb begin
end
endmodule
