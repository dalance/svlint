module noPrefix; // Module identifier of declaration should have prefix.
endmodule
