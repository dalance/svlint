module M;
  typedef enum int {
    i
  } E;
endmodule
