module A;
genvar i;
for(i=0;i<10;i++) begin
end
endmodule
