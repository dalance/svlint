module A;
Foo #() u_foo (a, b, c);
endmodule
