module M;
  initial begin
    unique0 case (a)
      default: b = 1;
    endcase
  end
endmodule
