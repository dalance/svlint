module A;
typedef enum logic {
    C
} B;
endmodule
