module M;
  always @(posedge clk) z--;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  always @(posedge clk) z++;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  always @* z = x + y--;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  always @* z = x + y++;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  genvar i;
  for (i = 4; i >= 0; i--) begin
    assign z[i] = y[i] + x[i];
  end
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  genvar i;
  for (i = 0; i < 5; i++) begin
    assign z[i] = y[i] + x[i];
  end
endmodule
