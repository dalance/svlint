module M (
  input
  a, // newline, not a space
  input    b, // too many spaces
  input/* comment */ c  // not a space
);
endmodule
