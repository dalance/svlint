module M;
	logic a;
endmodule
