module Bar;
endmodule