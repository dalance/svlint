class C;
  int Mn3; // Identifier doesn't match default required regex (lowercase).
endclass
