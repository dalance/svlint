module M;

logic [31:0] a;

endmodule
////////////////////////////////////////////////////////////////////////////////
module M;

logic [7:0][3:0] b;

endmodule
