program Bar;
endprogram