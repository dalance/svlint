module syntaxrules();
endmodule 


// Allowing Whitespace in Module Names
module syntaxrules ();
endmodule

// This testcase, when executed, is called from a file named "syntaxrules.module_identifier_matches_filename.pass.1of1"
// The rule matches all valid characters up until the first non-identifier (in this case, the period).
// The file identifier to be matched in this case becomes "syntaxrules" which matches the module identifier