module Xfoo; // Identifier doesn't match default forbidden regex (X prefix).
endmodule
