`default_nettype none
module M;
endmodule
