module A;
always_comb begin
end
always @ ( posedge a ) begin
end
endmodule
