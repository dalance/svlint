checker Xfoo; // Identifier doesn't match default forbidden regex (X prefix).
endchecker
