module M
  ( input  a
  , output b
  );
endmodule
