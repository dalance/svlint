module A(
    a,
    b
);
input  a;
output b;
endmodule
