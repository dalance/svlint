package Mn3; // Identifier doesn't match default required regex (lowercase).
endpackage
