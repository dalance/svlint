module A();
initial begin
    case (a)
        default: b = 1;
    endcase
end
endmodule
