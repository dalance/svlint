module M
  #( MN3 // Identifier matches default required regex (uppercase).
  ) ();
endmodule
