module A;
for(genvar i=0; i<10; i++) begin
end
endmodule
