package FooBar; endpackage
