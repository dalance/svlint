module A;
  function foo();
    if (a)
      return  ; // multiple spaces after `return`.
  endfunction
endmodule

