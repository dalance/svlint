package A;
parameter A = 1;
endpackage
