module A (
    inout tri a
);
endmodule
