module M;
  localparam L = 0;
endmodule
