module        M;
// End of line ^
endmodule
