module MN3 // Identifier matches default required regex (uppercase).
  ( a
  );
  input a;
endmodule
