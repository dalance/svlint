package P;
  localparam int A = 1;
endpackage
