module M;
  always_comb begin
  end
  always @(posedge a) begin
  end
endmodule
