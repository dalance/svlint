module A;
  always_comb
    case (x)
      1: a = 0;
    endcase
endmodule
