checker foo; // Unconfigured forbidden regex matches (almost) anything.
endchecker
