module M;
  A #(
  ) Mn3 (); // Identifier doesn't match default required regex (lowercase).
endmodule
