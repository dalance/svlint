module M;
  always @*
    assign c = a + b;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  always_comb
    assign c = a + b;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  always_latch
    assign c = a + b;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  always_ff @(posedge clk)
    assign c = a + b;
endmodule
