class foo; // Unconfigured forbidden regex matches (almost) anything.
endclass
