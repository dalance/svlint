module A;
function automatic A;
endfunction
endmodule
