package syntaxrules_package_identifier_matches_filename_pass_1of1;
endpackage

