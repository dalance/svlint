module A;
endmodule  : A // spaces immediately after `endmodule`
////////////////////////////////////////////////////////////////////////////////
package A;
endpackage  // multiple spaces then comment after `endpackage`
////////////////////////////////////////////////////////////////////////////////
interface A;
endinterface interface B; // space instead of newline after `endinterface`
endinterface
