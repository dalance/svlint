module M;
  Foo #() foo (a, b, c);
endmodule
