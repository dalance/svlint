module M;
  initial
    case (a)
      default: b = 1;
    endcase
endmodule
