interface foo; // Unconfigured forbidden regex matches (almost) anything.
endinterface
