module A;
wire a;
reg b;
endmodule
