`default_nettype none
module M;
endmodule
`default_nettype wire
