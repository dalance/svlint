module A #(parameter int a = 0) ();
endmodule
