program foo; // Unconfigured forbidden regex matches (almost) anything.
endprogram
