module mod_withPrefix; endmodule
