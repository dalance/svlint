module A;
function clog2;
endfunction
endmodule
