module M
  ( input var i_foo
  , input var logic [FOO-1:0] i_bar
  );
endmodule
