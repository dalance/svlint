module mN3; // Identifier matches default required regex (mixed-case).
endmodule
