module M;
  I #() u_foo (a, b, c);
endmodule
