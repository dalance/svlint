module M;
  function my_clog2;
  endfunction
endmodule
