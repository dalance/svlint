package P;
  localparam foo = 0; // Unconfigured forbidden regex matches (almost) anything.
endpackage
