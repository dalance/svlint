package fooBar; endpackage
