interface FooBar;
endinterface
