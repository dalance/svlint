module FooBar; endmodule
