module A (
    inout var a
);
endmodule
