module A (
    output var a
);
endmodule
