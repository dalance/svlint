class Xfoo; // Identifier doesn't match default forbidden regex (X prefix).
endclass
