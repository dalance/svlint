module A (
    test_if a,
    interface b
);
endmodule
