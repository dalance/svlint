module A
  #(parameter integer A = 32'b0
  ) ();
endmodule
////////////////////////////////////////////////////////////////////////////////
module A
  #(parameter logic B = 1'b0
  ) ();
endmodule
////////////////////////////////////////////////////////////////////////////////
module A
  #(parameter reg C = 1'b0
  , logic         Z = 1'b0 // TODO: Z isn't caught.
  ) ();
endmodule
