module M;
endmodule
