module M
  ( ref foo // Unconfigured forbidden regex matches (almost) anything.
  );
endmodule
