interface noPrefix;
endinterface
