module Mnonansi
  ( a
  , b
  );
  input  a;
  output b;
endmodule
