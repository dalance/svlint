interface Bar;
endinterface