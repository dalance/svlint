module A;
endmodule

