package pkg_withPrefix; endpackage
