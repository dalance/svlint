module A;
function A;
endfunction
endmodule
