module M;
  always_ff @(posedge clk)
    d <= q;
endmodule
