module A;
initial begin
for(int i=0;i<10;i++) begin
end
end
endmodule
