module M;

logic a [7:0];

endmodule;
////////////////////////////////////////////////////////////////////////////////
module M;

logic [31:0] b [0:7];

endmodule;
////////////////////////////////////////////////////////////////////////////////
module M;

localparam bit [7:0] ARRAY [0:3];

endmodule
////////////////////////////////////////////////////////////////////////////////
module M (
  input logic [7:0] a_in [0:5]
);

endmodule
