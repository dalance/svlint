module A();
  logic a;
endmodule
