module M;
  always @(a or b) q1 <= d;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  always_ff @(a, b or c) q2 <= d;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  always @( a
          or b
          , c
          ) q3 <= d;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  always_ff @(a
            , b
            or c
            ) q4 <= d;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  initial begin
    z = y;
    @(posedge a, negedge b, edge c or d)
    z = x;
  end
endmodule
