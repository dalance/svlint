module fooBar;
endmodule
