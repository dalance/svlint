module M;
  always_comb
    x <= 0;
endmodule
