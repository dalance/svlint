class C;
  function F;
    int mn3; // Identifier matches default required regex (lowercase).
  endfunction
endclass
