module A (
    inout wire a
);
endmodule
