module M
  ( a
  , b
  );
  input  a;
  output b;
endmodule
