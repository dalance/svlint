module M
  ( inout tri a
  );
endmodule
