module M;
  task foo; // Unconfigured forbidden regex matches (almost) anything.
  endtask
endmodule
