module aB3; // Identifier matches default required regex (mixed-case).
endmodule
