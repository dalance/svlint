module FooBar;
endmodule
