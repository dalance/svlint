module A();
initial begin
    unique case (a)
        default: b = 1;
    endcase
end
endmodule
