module M
  ( inout wire a
  );
endmodule
