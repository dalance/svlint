module A;
localparam a = 0;
endmodule
