module A;
always_ff if (x) y <= 0;
always_comb if (x) y = 0;
endmodule
