module A (
    input var a
);
endmodule
