module M;
  assign foo = bar    ; // Spaces preceeding semicolon.
endmodule
