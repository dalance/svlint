module M (
  input   a,
  inout   b   // multiple spaces after `input` or `inout` keywords
);
endmodule
