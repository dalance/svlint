class C;
  int foo; // Unconfigured forbidden regex matches (almost) anything.
endclass
