module M
  ( output var foo
  , output var logic [FOO-1:0] bar
  );
endmodule
