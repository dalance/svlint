interface I;
  modport mn3 // Identifier matches default required regex (lowercase).
  ( input i
  );
endinterface
