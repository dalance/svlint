module M;
  function F;
  endfunction
endmodule
