module A;
  Foo #() foo (a, b, c);
endmodule
