module M;
  task Mn3; // Identifier doesn't match default required regex (lowercase).
  endtask
endmodule
