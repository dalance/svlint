module M
  #(parameter a = 0
  ) ();
endmodule
////////////////////////////////////////////////////////////////////////////////
module M
  #(parameter a = int'(0)
  ) ();
endmodule
