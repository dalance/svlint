package P;
  function Mn3; // Identifier doesn't match default required regex (lowercase).
  endfunction
endpackage
