`default_nettype none
module A;
endmodule

