module M
  #( foo // Unconfigured forbidden regex matches (almost) anything.
  ) ();
endmodule
