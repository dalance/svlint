module foo; // Identifier matches default forbidden regex.
endmodule
