module A (
    input var i_a
);
endmodule
