module syntaxrules;
endmodule