package noPrefix; endpackage
