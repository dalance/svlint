module M;
  function clog2;
  endfunction
endmodule
