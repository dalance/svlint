module M;
  always @* a = b + c;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  always @(*) a = b + c;
endmodule
