module M;
  initial
    unique case (a)
      default: b = 1;
    endcase
endmodule
