interface noPrefix; endinterface
