class C;
  int Xfoo; // Identifier doesn't match default forbidden regex (X prefix).
endclass
