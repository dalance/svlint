module  A;
endmodule
