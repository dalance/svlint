module M
  ( output logic a
  );
endmodule
