module M
( inout var foo
, inout var logic [FOO-1:0] bar
);
endmodule
