module A;
always @* begin
end
always @ ( a or b ) begin
end
endmodule
