module foo; // Unconfigured forbidden regex matches (almost) anything.
endmodule
