module M
( output var o_foo
, output var logic [FOO-1:0] o_bar
);
endmodule
