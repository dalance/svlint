interface mn3; // Identifier matches default required regex (lowercase).
endinterface
