package P;
  parameter int A = 1;
endpackage
