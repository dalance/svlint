module M;
  always_comb z = x + y;
endmodule
