module mn3 // Identifier doesn't match default required regex (uppercase).
  ( a
  );
  input a;
endmodule
