package mn3; // Identifier matches default required regex (lowercase).
endpackage
