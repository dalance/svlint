module A;
generate
endgenerate
endmodule
