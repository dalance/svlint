module A (
    inout var b_a
);
endmodule
