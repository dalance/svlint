module fooBar; endmodule
