module noPrefix; endmodule
