module M
  #(parameter int P = 0
  ) ();
endmodule
