// Copyright (c) 1234 HOLDER
// The string "Copyright" is lowercase but capitalized.
// The symbol "(c)" may be either uppercase or lowercase.
////////////////////////////////////////////////////////////////////////////////
// copyright (c) 1234 HOLDER
// The string "copyright" is fully lowercase.
////////////////////////////////////////////////////////////////////////////////
// COPYRIGHT   (C)    1234    HOLDER
// The string "COPYRIGHT" is fully uppercase.
// Components may be separated by multiple spaces.
////////////////////////////////////////////////////////////////////////////////
// foo bar Copyright (c) 1234 HOLDER foo bar
// There may be other text on either end of the same line.
