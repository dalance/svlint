module M;
  if (a) begin
  end
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  case (a)
      default: a;
  endcase
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  for (genvar i=0; i < 10; i++) begin
  end
endmodule
