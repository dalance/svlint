/*
Lorem ipsum dolor sit amet, consectetur adipiscing elit, sed do eiusmod    GOOD><BAD
tempor incididunt ut labore et dolore magna aliqua. Ut enim ad minim veniam,
quis nostrud exercitation ullamco laboris nisi ut aliquip ex ea commodo    GOOD><BAD
consequat. Duis aute irure dolor in reprehenderit in voluptate velit esse  GOOD><BAD
Zażółć gęślą jaźń                                                          GOOD><BAD
foo                                                                        GOOD><BAD
cillum dolore eu fugiat nulla pariatur. Excepteur sint occaecat cupidatat non
proident, sunt in culpa qui officia deserunt mollit anim id est laborum.
*/
