module A;
logic a;
logic b;
endmodule
