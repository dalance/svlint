package FooBar;
endpackage
