package fooBar;
endpackage
