module M
  ( inout var b_foo
  , input var logic [FOO-1:0] b_bar
  );
endmodule
