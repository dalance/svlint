interface fooBar; endinterface
