program syntaxrules_program_identifier_matches_filename_pass_1of1;
endprogram