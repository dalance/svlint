module Ab3; // Identifier doesn't match default required regex (mixed-case).
endmodule
