module M
  #( Mn3 // Identifier doesn't match default required regex (uppercase).
  ) ();
endmodule
