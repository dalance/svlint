module A #(parameter a = 0) ();
endmodule
