package P;
  localparam MN3 = 0; // Identifier matches default required regex (uppercase).
endpackage
