module M;
  always @* begin
  end
endmodule
