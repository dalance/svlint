module A(
    input  a,
    output b
);
endmodule
