module M;
endmodule  : M // spaces immediately after `endmodule`
////////////////////////////////////////////////////////////////////////////////
package P;
endpackage  // multiple spaces then comment after `endpackage`
////////////////////////////////////////////////////////////////////////////////
interface I;
endinterface interface J; // space instead of newline after `endinterface`
endinterface
