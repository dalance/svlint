package A;
localparam A = 1;
endpackage
