program mn3; // Identifier matches default required regex (lowercase).
endprogram
