package M;
  localparam int A = 1;
endpackage
