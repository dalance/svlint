package foo; // Unconfigured forbidden regex matches (almost) anything.
endpackage
