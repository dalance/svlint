module A (
    input logic a
);
endmodule
