module M;
                
// End of line ^
endmodule

module M;       
// End of line ^
endmodule
