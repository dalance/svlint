module M;

logic a [7:0];

endmodule;
////////////////////////////////////////////////////////////////////////////////
module M;

logic [31:0] b [0:7];

endmodule;
