module syntaxrules_module_identifier_matches_filename_pass_1of1;
endmodule