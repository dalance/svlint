module M;
  always @(posedge clk) z = z - 1;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  always @(posedge clk) z = z + 1;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  always @* z = z - 1;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  always @* z = z + 1;
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  genvar i;
  for (i = 4; i >= 0; i = i - 1) begin
    assign z[i] = y[i] + x[i];
  end
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  genvar i;
  for (i = 0; i < 5; i = i + 1) begin
    assign z[i] = y[i] + x[i];
  end
endmodule
