module M;
  localparam int P1 = a | b; // Single space around `|`.

  localparam int P2 = a & aMask; // Single space before `&`.
endmodule
