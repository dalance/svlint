module M;
  task mn3; // Identifier matches default required regex (lowercase).
  endtask
endmodule
