`default_nettype none
module M;
endmodule
////////////////////////////////////////////////////////////////////////////////
/* svlint off default_nettype_none */
module M;
endmodule
/* svlint on default_nettype_none */
