module A;
always_comb begin
    x = 0;
end
endmodule
