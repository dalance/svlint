module M (
  input a,
  inout b,
  input  c,
  inout  d,
  output e
);
endmodule
