module A;
localparam int a = 0;
endmodule
