module M
  ( test_if a
  );
endmodule
////////////////////////////////////////////////////////////////////////////////
module M
  ( interface b
  );
endmodule
