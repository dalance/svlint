module M
  #(parameter int a = 0
  ) ();
endmodule
