localparam int A = 1;
