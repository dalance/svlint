module A (
    output var o_a
);
endmodule
