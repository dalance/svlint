package noPrefix;
endpackage
