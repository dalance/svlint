module M;
  typedef enum
    { i
    } E;
endmodule
