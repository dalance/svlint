program syntaxrules;
endprogram