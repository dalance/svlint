package syntaxrules;
endpackage

