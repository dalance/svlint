module M;
  always_comb begin
  end
endmodule
