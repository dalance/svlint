module M;
  initial
    for(int i=0; i < 10; i++) begin
    end
endmodule
