module M;
  generate
  endgenerate
endmodule
