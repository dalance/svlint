module M;
  assign foo = bar; // No space preceeding semicolon.
endmodule
