module M;
  localparam integer A = 32'b0; // 32b
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  localparam logic B = 1'b0; // 1b
endmodule
////////////////////////////////////////////////////////////////////////////////
module M;
  localparam reg C = 1'b0; // 1b
endmodule
