module A;
typedef enum {
    C
} B;
endmodule
