module M
  ( input var foo
  , input var logic [FOO-1:0] bar
  );
endmodule
