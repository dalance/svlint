module M;
  always @* z = x + y;
endmodule
