module Mansi
  ( input  a
  , output b
  );
endmodule

module Mansi_noPort;
endmodule

module Mansi_defaultInout
  ( a
  , b
  );
endmodule
