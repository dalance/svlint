interface syntaxrules;
endinterface