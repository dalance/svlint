module M;
  A #(
  ) foo (); // Unconfigured forbidden regex matches (almost) anything.
endmodule
