module A;
function my_clog2;
endfunction
endmodule
