module M;
  always @(posedge clk)
    d <= q;
endmodule
