interface syntaxrules_interface_identifier_matches_filename_pass_1of1;
endinterface