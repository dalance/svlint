package P;
  function mn3; // Identifier matches default required regex (lowercase).
  endfunction
endpackage
