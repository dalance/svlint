module M;
  localparam int A = 0;
endmodule
