module M
  ( output var logic a
  );
endmodule
