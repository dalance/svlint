module M
  ( input logic a
  );
endmodule
