module A (
    output logic a
);
endmodule
