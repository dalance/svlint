module A (
    test_if.a a,
    interface.b b
);
endmodule
