checker mn3; // Identifier matches default required regex (lowercase).
endchecker
