interface ifc_withPrefix;
endinterface
