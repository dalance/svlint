package P;
  function foo; // Unconfigured forbidden regex matches (almost) anything.
  endfunction
endpackage
