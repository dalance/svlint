module A;
always_ff begin
    x = 0;
end
endmodule
