module M;
  wire a;
  reg b;
endmodule
