interface fooBar;
endinterface
