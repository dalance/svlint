module A;
endmodule
