module foo // Unconfigured forbidden regex matches (almost) anything.
  ( a
  );
  input a;
endmodule
