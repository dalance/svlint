package P;
  localparam Mn3 = 0; // Identifier doesn't match default required regex (uppercase).
endpackage
