module M;
  A #(
  ) mn3 (); // Identifier matches default required regex (lowercase).
endmodule
