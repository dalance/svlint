module M;
  for (genvar i=0; i < 10; i++) begin: l_foo
  end: l_foo
endmodule
