module A;
if (a) begin
end else if (a) begin
end else begin
end
endmodule
