module M;
  initial begin
    int i;
    for(i=0; i < 10; i++) begin
    end
  end
endmodule
