interface FooBar; endinterface
