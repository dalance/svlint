module A;
if (a) begin: a
end else if (b) begin: a
end else begin: a
end
endmodule
