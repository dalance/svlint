module M;
  for(genvar i=0; i < 10; i++) begin: a
  end
endmodule
