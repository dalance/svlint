package P;
  localparam int A = 1;
endpackage
////////////////////////////////////////////////////////////////////////////////
package foo;
   class bar #( parameter int baz );
   endclass
endpackage
