module M
  ( input var a
  );
endmodule
